package pkg_strings;
    parameter S_CRLF = 9'd0;
    parameter S_hello_world = 9'd3;
    parameter S_startup_message = 9'd16;
    parameter S_waiting = 9'd46;
    parameter S_detect_full = 9'd72;
    parameter S_detect_low = 9'd100;
endpackage
