package pkg_strings;
    parameter S_hello_world = 9'd0;
    parameter S_startup_message = 9'd13;
endpackage
