
module strings(
    input               clk,
    input               rd,
    input       [8:0]   raddr,
    input               wr,
    input       [8:0]   waddr,
    input       [7:0]   din,
    output reg  [7:0]   dout
);

    reg [7:0] ram [511:0];

    always @(posedge clk) begin
        if (rd)
            dout <= ram[raddr];
        if (wr)
            ram[waddr] <= din;
    end

    initial begin
        ram[0] = 8'd72; // H
        ram[1] = 8'd101; // e
        ram[2] = 8'd108; // l
        ram[3] = 8'd108; // l
        ram[4] = 8'd111; // o
        ram[5] = 8'd32; //  
        ram[6] = 8'd119; // w
        ram[7] = 8'd111; // o
        ram[8] = 8'd114; // r
        ram[9] = 8'd108; // l
        ram[10] = 8'd100; // d
        ram[11] = 8'd33; // !
        ram[12] = 8'd0;
        ram[13] = 8'd126; // ~
        ram[14] = 8'd126; // ~
        ram[15] = 8'd126; // ~
        ram[16] = 8'd87; // W
        ram[17] = 8'd101; // e
        ram[18] = 8'd108; // l
        ram[19] = 8'd99; // c
        ram[20] = 8'd111; // o
        ram[21] = 8'd109; // m
        ram[22] = 8'd101; // e
        ram[23] = 8'd32; //  
        ram[24] = 8'd116; // t
        ram[25] = 8'd111; // o
        ram[26] = 8'd32; //  
        ram[27] = 8'd83; // S
        ram[28] = 8'd108; // l
        ram[29] = 8'd111; // o
        ram[30] = 8'd119; // w
        ram[31] = 8'd119; // w
        ram[32] = 8'd111; // o
        ram[33] = 8'd114; // r
        ram[34] = 8'd109; // m
        ram[35] = 8'd32; //  
        ram[36] = 8'd85; // U
        ram[37] = 8'd83; // S
        ram[38] = 8'd66; // B
        ram[39] = 8'd126; // ~
        ram[40] = 8'd126; // ~
        ram[41] = 8'd126; // ~
        ram[42] = 8'd0;
        ram[43] = 8'd0;
        ram[44] = 8'd0;
        ram[45] = 8'd0;
        ram[46] = 8'd0;
        ram[47] = 8'd0;
        ram[48] = 8'd0;
        ram[49] = 8'd0;
        ram[50] = 8'd0;
        ram[51] = 8'd0;
        ram[52] = 8'd0;
        ram[53] = 8'd0;
        ram[54] = 8'd0;
        ram[55] = 8'd0;
        ram[56] = 8'd0;
        ram[57] = 8'd0;
        ram[58] = 8'd0;
        ram[59] = 8'd0;
        ram[60] = 8'd0;
        ram[61] = 8'd0;
        ram[62] = 8'd0;
        ram[63] = 8'd0;
        ram[64] = 8'd0;
        ram[65] = 8'd0;
        ram[66] = 8'd0;
        ram[67] = 8'd0;
        ram[68] = 8'd0;
        ram[69] = 8'd0;
        ram[70] = 8'd0;
        ram[71] = 8'd0;
        ram[72] = 8'd0;
        ram[73] = 8'd0;
        ram[74] = 8'd0;
        ram[75] = 8'd0;
        ram[76] = 8'd0;
        ram[77] = 8'd0;
        ram[78] = 8'd0;
        ram[79] = 8'd0;
        ram[80] = 8'd0;
        ram[81] = 8'd0;
        ram[82] = 8'd0;
        ram[83] = 8'd0;
        ram[84] = 8'd0;
        ram[85] = 8'd0;
        ram[86] = 8'd0;
        ram[87] = 8'd0;
        ram[88] = 8'd0;
        ram[89] = 8'd0;
        ram[90] = 8'd0;
        ram[91] = 8'd0;
        ram[92] = 8'd0;
        ram[93] = 8'd0;
        ram[94] = 8'd0;
        ram[95] = 8'd0;
        ram[96] = 8'd0;
        ram[97] = 8'd0;
        ram[98] = 8'd0;
        ram[99] = 8'd0;
        ram[100] = 8'd0;
        ram[101] = 8'd0;
        ram[102] = 8'd0;
        ram[103] = 8'd0;
        ram[104] = 8'd0;
        ram[105] = 8'd0;
        ram[106] = 8'd0;
        ram[107] = 8'd0;
        ram[108] = 8'd0;
        ram[109] = 8'd0;
        ram[110] = 8'd0;
        ram[111] = 8'd0;
        ram[112] = 8'd0;
        ram[113] = 8'd0;
        ram[114] = 8'd0;
        ram[115] = 8'd0;
        ram[116] = 8'd0;
        ram[117] = 8'd0;
        ram[118] = 8'd0;
        ram[119] = 8'd0;
        ram[120] = 8'd0;
        ram[121] = 8'd0;
        ram[122] = 8'd0;
        ram[123] = 8'd0;
        ram[124] = 8'd0;
        ram[125] = 8'd0;
        ram[126] = 8'd0;
        ram[127] = 8'd0;
        ram[128] = 8'd0;
        ram[129] = 8'd0;
        ram[130] = 8'd0;
        ram[131] = 8'd0;
        ram[132] = 8'd0;
        ram[133] = 8'd0;
        ram[134] = 8'd0;
        ram[135] = 8'd0;
        ram[136] = 8'd0;
        ram[137] = 8'd0;
        ram[138] = 8'd0;
        ram[139] = 8'd0;
        ram[140] = 8'd0;
        ram[141] = 8'd0;
        ram[142] = 8'd0;
        ram[143] = 8'd0;
        ram[144] = 8'd0;
        ram[145] = 8'd0;
        ram[146] = 8'd0;
        ram[147] = 8'd0;
        ram[148] = 8'd0;
        ram[149] = 8'd0;
        ram[150] = 8'd0;
        ram[151] = 8'd0;
        ram[152] = 8'd0;
        ram[153] = 8'd0;
        ram[154] = 8'd0;
        ram[155] = 8'd0;
        ram[156] = 8'd0;
        ram[157] = 8'd0;
        ram[158] = 8'd0;
        ram[159] = 8'd0;
        ram[160] = 8'd0;
        ram[161] = 8'd0;
        ram[162] = 8'd0;
        ram[163] = 8'd0;
        ram[164] = 8'd0;
        ram[165] = 8'd0;
        ram[166] = 8'd0;
        ram[167] = 8'd0;
        ram[168] = 8'd0;
        ram[169] = 8'd0;
        ram[170] = 8'd0;
        ram[171] = 8'd0;
        ram[172] = 8'd0;
        ram[173] = 8'd0;
        ram[174] = 8'd0;
        ram[175] = 8'd0;
        ram[176] = 8'd0;
        ram[177] = 8'd0;
        ram[178] = 8'd0;
        ram[179] = 8'd0;
        ram[180] = 8'd0;
        ram[181] = 8'd0;
        ram[182] = 8'd0;
        ram[183] = 8'd0;
        ram[184] = 8'd0;
        ram[185] = 8'd0;
        ram[186] = 8'd0;
        ram[187] = 8'd0;
        ram[188] = 8'd0;
        ram[189] = 8'd0;
        ram[190] = 8'd0;
        ram[191] = 8'd0;
        ram[192] = 8'd0;
        ram[193] = 8'd0;
        ram[194] = 8'd0;
        ram[195] = 8'd0;
        ram[196] = 8'd0;
        ram[197] = 8'd0;
        ram[198] = 8'd0;
        ram[199] = 8'd0;
        ram[200] = 8'd0;
        ram[201] = 8'd0;
        ram[202] = 8'd0;
        ram[203] = 8'd0;
        ram[204] = 8'd0;
        ram[205] = 8'd0;
        ram[206] = 8'd0;
        ram[207] = 8'd0;
        ram[208] = 8'd0;
        ram[209] = 8'd0;
        ram[210] = 8'd0;
        ram[211] = 8'd0;
        ram[212] = 8'd0;
        ram[213] = 8'd0;
        ram[214] = 8'd0;
        ram[215] = 8'd0;
        ram[216] = 8'd0;
        ram[217] = 8'd0;
        ram[218] = 8'd0;
        ram[219] = 8'd0;
        ram[220] = 8'd0;
        ram[221] = 8'd0;
        ram[222] = 8'd0;
        ram[223] = 8'd0;
        ram[224] = 8'd0;
        ram[225] = 8'd0;
        ram[226] = 8'd0;
        ram[227] = 8'd0;
        ram[228] = 8'd0;
        ram[229] = 8'd0;
        ram[230] = 8'd0;
        ram[231] = 8'd0;
        ram[232] = 8'd0;
        ram[233] = 8'd0;
        ram[234] = 8'd0;
        ram[235] = 8'd0;
        ram[236] = 8'd0;
        ram[237] = 8'd0;
        ram[238] = 8'd0;
        ram[239] = 8'd0;
        ram[240] = 8'd0;
        ram[241] = 8'd0;
        ram[242] = 8'd0;
        ram[243] = 8'd0;
        ram[244] = 8'd0;
        ram[245] = 8'd0;
        ram[246] = 8'd0;
        ram[247] = 8'd0;
        ram[248] = 8'd0;
        ram[249] = 8'd0;
        ram[250] = 8'd0;
        ram[251] = 8'd0;
        ram[252] = 8'd0;
        ram[253] = 8'd0;
        ram[254] = 8'd0;
        ram[255] = 8'd0;
        ram[256] = 8'd0;
        ram[257] = 8'd0;
        ram[258] = 8'd0;
        ram[259] = 8'd0;
        ram[260] = 8'd0;
        ram[261] = 8'd0;
        ram[262] = 8'd0;
        ram[263] = 8'd0;
        ram[264] = 8'd0;
        ram[265] = 8'd0;
        ram[266] = 8'd0;
        ram[267] = 8'd0;
        ram[268] = 8'd0;
        ram[269] = 8'd0;
        ram[270] = 8'd0;
        ram[271] = 8'd0;
        ram[272] = 8'd0;
        ram[273] = 8'd0;
        ram[274] = 8'd0;
        ram[275] = 8'd0;
        ram[276] = 8'd0;
        ram[277] = 8'd0;
        ram[278] = 8'd0;
        ram[279] = 8'd0;
        ram[280] = 8'd0;
        ram[281] = 8'd0;
        ram[282] = 8'd0;
        ram[283] = 8'd0;
        ram[284] = 8'd0;
        ram[285] = 8'd0;
        ram[286] = 8'd0;
        ram[287] = 8'd0;
        ram[288] = 8'd0;
        ram[289] = 8'd0;
        ram[290] = 8'd0;
        ram[291] = 8'd0;
        ram[292] = 8'd0;
        ram[293] = 8'd0;
        ram[294] = 8'd0;
        ram[295] = 8'd0;
        ram[296] = 8'd0;
        ram[297] = 8'd0;
        ram[298] = 8'd0;
        ram[299] = 8'd0;
        ram[300] = 8'd0;
        ram[301] = 8'd0;
        ram[302] = 8'd0;
        ram[303] = 8'd0;
        ram[304] = 8'd0;
        ram[305] = 8'd0;
        ram[306] = 8'd0;
        ram[307] = 8'd0;
        ram[308] = 8'd0;
        ram[309] = 8'd0;
        ram[310] = 8'd0;
        ram[311] = 8'd0;
        ram[312] = 8'd0;
        ram[313] = 8'd0;
        ram[314] = 8'd0;
        ram[315] = 8'd0;
        ram[316] = 8'd0;
        ram[317] = 8'd0;
        ram[318] = 8'd0;
        ram[319] = 8'd0;
        ram[320] = 8'd0;
        ram[321] = 8'd0;
        ram[322] = 8'd0;
        ram[323] = 8'd0;
        ram[324] = 8'd0;
        ram[325] = 8'd0;
        ram[326] = 8'd0;
        ram[327] = 8'd0;
        ram[328] = 8'd0;
        ram[329] = 8'd0;
        ram[330] = 8'd0;
        ram[331] = 8'd0;
        ram[332] = 8'd0;
        ram[333] = 8'd0;
        ram[334] = 8'd0;
        ram[335] = 8'd0;
        ram[336] = 8'd0;
        ram[337] = 8'd0;
        ram[338] = 8'd0;
        ram[339] = 8'd0;
        ram[340] = 8'd0;
        ram[341] = 8'd0;
        ram[342] = 8'd0;
        ram[343] = 8'd0;
        ram[344] = 8'd0;
        ram[345] = 8'd0;
        ram[346] = 8'd0;
        ram[347] = 8'd0;
        ram[348] = 8'd0;
        ram[349] = 8'd0;
        ram[350] = 8'd0;
        ram[351] = 8'd0;
        ram[352] = 8'd0;
        ram[353] = 8'd0;
        ram[354] = 8'd0;
        ram[355] = 8'd0;
        ram[356] = 8'd0;
        ram[357] = 8'd0;
        ram[358] = 8'd0;
        ram[359] = 8'd0;
        ram[360] = 8'd0;
        ram[361] = 8'd0;
        ram[362] = 8'd0;
        ram[363] = 8'd0;
        ram[364] = 8'd0;
        ram[365] = 8'd0;
        ram[366] = 8'd0;
        ram[367] = 8'd0;
        ram[368] = 8'd0;
        ram[369] = 8'd0;
        ram[370] = 8'd0;
        ram[371] = 8'd0;
        ram[372] = 8'd0;
        ram[373] = 8'd0;
        ram[374] = 8'd0;
        ram[375] = 8'd0;
        ram[376] = 8'd0;
        ram[377] = 8'd0;
        ram[378] = 8'd0;
        ram[379] = 8'd0;
        ram[380] = 8'd0;
        ram[381] = 8'd0;
        ram[382] = 8'd0;
        ram[383] = 8'd0;
        ram[384] = 8'd0;
        ram[385] = 8'd0;
        ram[386] = 8'd0;
        ram[387] = 8'd0;
        ram[388] = 8'd0;
        ram[389] = 8'd0;
        ram[390] = 8'd0;
        ram[391] = 8'd0;
        ram[392] = 8'd0;
        ram[393] = 8'd0;
        ram[394] = 8'd0;
        ram[395] = 8'd0;
        ram[396] = 8'd0;
        ram[397] = 8'd0;
        ram[398] = 8'd0;
        ram[399] = 8'd0;
        ram[400] = 8'd0;
        ram[401] = 8'd0;
        ram[402] = 8'd0;
        ram[403] = 8'd0;
        ram[404] = 8'd0;
        ram[405] = 8'd0;
        ram[406] = 8'd0;
        ram[407] = 8'd0;
        ram[408] = 8'd0;
        ram[409] = 8'd0;
        ram[410] = 8'd0;
        ram[411] = 8'd0;
        ram[412] = 8'd0;
        ram[413] = 8'd0;
        ram[414] = 8'd0;
        ram[415] = 8'd0;
        ram[416] = 8'd0;
        ram[417] = 8'd0;
        ram[418] = 8'd0;
        ram[419] = 8'd0;
        ram[420] = 8'd0;
        ram[421] = 8'd0;
        ram[422] = 8'd0;
        ram[423] = 8'd0;
        ram[424] = 8'd0;
        ram[425] = 8'd0;
        ram[426] = 8'd0;
        ram[427] = 8'd0;
        ram[428] = 8'd0;
        ram[429] = 8'd0;
        ram[430] = 8'd0;
        ram[431] = 8'd0;
        ram[432] = 8'd0;
        ram[433] = 8'd0;
        ram[434] = 8'd0;
        ram[435] = 8'd0;
        ram[436] = 8'd0;
        ram[437] = 8'd0;
        ram[438] = 8'd0;
        ram[439] = 8'd0;
        ram[440] = 8'd0;
        ram[441] = 8'd0;
        ram[442] = 8'd0;
        ram[443] = 8'd0;
        ram[444] = 8'd0;
        ram[445] = 8'd0;
        ram[446] = 8'd0;
        ram[447] = 8'd0;
        ram[448] = 8'd0;
        ram[449] = 8'd0;
        ram[450] = 8'd0;
        ram[451] = 8'd0;
        ram[452] = 8'd0;
        ram[453] = 8'd0;
        ram[454] = 8'd0;
        ram[455] = 8'd0;
        ram[456] = 8'd0;
        ram[457] = 8'd0;
        ram[458] = 8'd0;
        ram[459] = 8'd0;
        ram[460] = 8'd0;
        ram[461] = 8'd0;
        ram[462] = 8'd0;
        ram[463] = 8'd0;
        ram[464] = 8'd0;
        ram[465] = 8'd0;
        ram[466] = 8'd0;
        ram[467] = 8'd0;
        ram[468] = 8'd0;
        ram[469] = 8'd0;
        ram[470] = 8'd0;
        ram[471] = 8'd0;
        ram[472] = 8'd0;
        ram[473] = 8'd0;
        ram[474] = 8'd0;
        ram[475] = 8'd0;
        ram[476] = 8'd0;
        ram[477] = 8'd0;
        ram[478] = 8'd0;
        ram[479] = 8'd0;
        ram[480] = 8'd0;
        ram[481] = 8'd0;
        ram[482] = 8'd0;
        ram[483] = 8'd0;
        ram[484] = 8'd0;
        ram[485] = 8'd0;
        ram[486] = 8'd0;
        ram[487] = 8'd0;
        ram[488] = 8'd0;
        ram[489] = 8'd0;
        ram[490] = 8'd0;
        ram[491] = 8'd0;
        ram[492] = 8'd0;
        ram[493] = 8'd0;
        ram[494] = 8'd0;
        ram[495] = 8'd0;
        ram[496] = 8'd0;
        ram[497] = 8'd0;
        ram[498] = 8'd0;
        ram[499] = 8'd0;
        ram[500] = 8'd0;
        ram[501] = 8'd0;
        ram[502] = 8'd0;
        ram[503] = 8'd0;
        ram[504] = 8'd0;
        ram[505] = 8'd0;
        ram[506] = 8'd0;
        ram[507] = 8'd0;
        ram[508] = 8'd0;
        ram[509] = 8'd0;
        ram[510] = 8'd0;
        ram[511] = 8'd0;
    end
endmodule
